interface intf_rst ();
	bit rst_in;
	bit rst_out;
endinterface : intf_rst