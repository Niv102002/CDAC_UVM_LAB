class agent_master extends uvm_agent;

`uvm_component_utlis(agent_master)

monitor_master mon_m;
sequencer_master seqr_m;

endclass : agent_master